// This file contains multiple modules that will have to be used a lot, such as a register, multiplexer, multiplier, adder, comparator, etc.